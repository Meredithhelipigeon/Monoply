0
0 0 0 0 0 r h 0 B 17 B 
0 0 0 0 0 r h 4 B 10 B 


2 2 1 5 4 6 1 3 2 3 0 3 3 3 0 4 2 4 1 11 4 11 0 8 0 8 3 11 3 8 1 11 4 9 5 7 2 12 
-1
